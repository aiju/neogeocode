`default_nettype none
`define CLKMUL 8
`define CLKDIV 5
`define MHZ (100.0*`CLKMUL/`CLKDIV)
